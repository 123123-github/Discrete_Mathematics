/*
    date:   2018/06/02
    tag:    test sl2
*/

module t_sl2();
    reg[31:0]   a;
    reg[25:0]   b;

    wire[31:0]  m;
    wire[25:0]  n;

    initial
    fork
        #50 a = 32'h8fff0000;   // 1000_1111_1111_1111_0000...0000  -> 3ffc0000
        #50 b = 26'h83000000;   // 1000_00,11_0000...0000
        
        #150 a = 32'hff002222;
        #150 b = 26'h55555555;
        
        #250 a = 32'h5f012222;
        #250 b = 26'h66666666;        
        
    join

    sl2 #(32) SL2_32( .a(a), .y(m));
    sl2 #(26) SL2_26( .a(b), .y(n));


endmodule